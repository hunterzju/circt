module ALU();
endmodule
